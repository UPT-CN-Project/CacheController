//==============================================================================
// Module: bitwise_comparator
// Description:
//   Compares two multi-bit vectors, `in_0` and `in_1`, and outputs `eq` which
//   is high (1) if and only if all corresponding bits in the two vectors match.
//   Internally, it instantiates a `bit_comparator` for each bit position to
//   produce a per-bit equality vector `bitwise_eq`. That vector is then fed to
//   an `and_wordgate` to ensure every bit comparison is true.
//
// Parameters:
//   w  - Width of the input vectors `in_0` and `in_1`. Determines how many
//        bits get compared. Default is 8.
//
// Ports:
//   input  [w-1:0] in_0
//     - First multi-bit input vector to compare.
//   input  [w-1:0] in_1
//     - Second multi-bit input vector to compare.
//   output        eq
//     - Single-bit output: high if in_0 == in_1 on every bit, low otherwise.
//
// Internal Signals:
//   wire [w-1:0] bitwise_eq
//     - A bus of per-bit equality results. bitwise_eq[i] is 1 if in_0[i] == in_1[i],
//       0 otherwise. This bus is generated by instantiating `w` copies of
//       `bit_comparator`.
//
// Behavior:
//   1. For each bit index i from 0 to w-1:
//        bitwise_eq[i] = 1 if in_0[i] == in_1[i], else 0.
//   2. The `and_wordgate` reduction ANDs all bits of `bitwise_eq`. If every bit
//      matches (all bitwise_eq bits are 1), then `eq` = 1. If any bit differs,
//      `eq` = 0.
//
// Usage Notes:
//   - Use this module when you need a vector-wide equality check in purely
//     structural form (instantiating bitwise comparators and a reduction AND).
//   - Synthesizable and parameterizable to any width.
//
// Example Instantiation (for 16-bit comparison):
//   bitwise_comparator #(.w(16)) u_bcmp (
//       .in_0 (data_from_cache),
//       .in_1 (address_tag),
//       .eq   (tags_match_signal)
//   );
//
//==============================================================================

module bitwise_comparator #(
    parameter w = 8  // Width of input vectors
) (
    input  wire [w-1:0] in_0,  // First input vector
    input  wire [w-1:0] in_1,  // Second input vector
    output              eq     // High if all bits match
);

    // A vector of per-bit equality results.
    // bitwise_eq[i] == 1 if in_0[i] == in_1[i], else 0.
    wire [w-1:0] bitwise_eq;

    // Generate block: instantiate a `bit_comparator` for each bit position
    // from 0..w-1, wiring in_0[i], in_1[i] into eq[i].
    generate
        genvar i;
        for (i = 0; i < w; i = i + 1) begin : comp_instances
            bit_comparator uut (
                .b0(in_0[i]),
                .b1(in_1[i]),
                .eq(bitwise_eq[i])
            );
        end
    endgenerate

    // Reduction AND: if every bitwise_eq[i] is 1, then eq = 1. Otherwise 0.
    and_wordgate #(
        .w(w)
    ) reduction_and (
        .in  (bitwise_eq),
        .AND_(eq)
    );

endmodule
