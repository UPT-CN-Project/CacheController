// The four_way_set module implements a four-way set associative cache set.
// It manages multiple cache lines within a set, handles read and write operations, updates cache line ages, and determines cache hits or misses.
// Four instances of the cache_line module handle the actual data storage and retrieval.
// Each cache line operates based on the provided signals (try_read, try_write, reset_age, increment_age).
// The mux4to1 modules select the appropriate data and hit/miss signals based on the sel signal generated by the encoder4to2 module.
// The hit_miss_set output is directly assigned from line_hit_miss.

module four_way_set #(
    parameter ADDRESS_WORD_SIZE = 32,
    parameter TAG_SIZE          = 19,
    parameter BLOCK_SIZE        = 16,
    parameter WORD_SIZE         = 4
) (
    input wire                         clk,
    input wire                         rst_b,
    input wire [ADDRESS_WORD_SIZE-1:0] address_word,
    input wire                         try_read,
    input wire                         try_write,
    input wire [                  7:0] write_data,
    input wire [                  3:0] reset_age,     // per‐way “reset age” pulses
    input wire [                  3:0] increment_age, // per‐way “increment age” pulses

    output wire [7:0] data,         // selected byte from the chosen way
    output wire [7:0] ages,         // concatenated {way3_age, way2_age, way1_age, way0_age}
    output wire       hit_miss,     // 1 if the chosen way hits
    output wire [3:0] hit_miss_set  // one‐hot of which way(s) hit
);

    //----------------------------------------------------------------------
    // Internal “select” register (one-hot).  Each bit = “give this way the next
    // operation (read/write) permission.”
    //----------------------------------------------------------------------
    reg  [ 3:0] ready;

    //----------------------------------------------------------------------
    // Collate all 4 lines’ data, hit/miss, empty, age signals into buses:
    //----------------------------------------------------------------------
    wire [31:0] line_data;  // 4 × 8‐bit “data out” buses concatenated
    wire [ 3:0] line_hit_miss;  // each way’s hit/miss flag (1 = this way hit)
    wire [ 3:0] line_is_empty;  // each way’s “empty?” flag (1 = line is not valid)
    wire [ 1:0] sel;  // 2‐bit index = which bit of “ready” is set

    //----------------------------------------------------------------------
    // 4‐to‐2 encoder: if ready=4'b0100, then sel=2'b10.  If ready=4'b0000,
    // we define sel=2'b00 (default to way0).
    //----------------------------------------------------------------------
    encoder4to2 enc4to2_inst (
        .in (ready),
        .out(sel)
    );

    //----------------------------------------------------------------------
    // Instantiate four cache_line modules.  Each way sees:
    //   - clk, rst_b, its own “ready[i]” bit, the global address_word,
    //   - the global try_read/try_write/write_data signals,
    //   - reset_age[i] and increment_age[i],
    //   - and returns an 8‐bit “data” slice, 2‐bit “age,” 1‐bit “hit_miss,”
    //     and 1‐bit “is_empty.”
    //----------------------------------------------------------------------
    generate
        genvar i;
        for (i = 0; i < 4; i = i + 1) begin : cache_lines
            cache_line #(
                .ADDRESS_WORD_SIZE(ADDRESS_WORD_SIZE),
                .TAG_SIZE         (TAG_SIZE),
                .BLOCK_SIZE       (BLOCK_SIZE),
                .WORD_SIZE        (WORD_SIZE)
            ) line_inst (
                .clk          (clk),
                .rst_b        (rst_b),
                .ready        (ready[i]),
                .address_word (address_word),
                .try_read     (try_read),
                .try_write    (try_write),
                .write_data   (write_data),
                .reset_age    (reset_age[i]),
                .increment_age(increment_age[i]),

                .data    (line_data[8*(i+1)-1 : 8*i]),  // way i → bits [8*i +: 8]
                .age     (ages[2*i+1 : 2*i]),           // way i → bits [2*i +: 2]
                .hit_miss(line_hit_miss[i]),
                .is_empty(line_is_empty[i])
            );
        end
    endgenerate

    //----------------------------------------------------------------------
    // Convey “which way hit” as a one‐hot vector.  If multiple ways somehow
    // flagged a hit simultaneously (shouldn’t happen in a correct cache),
    // then hit_miss_set will show them all.
    //----------------------------------------------------------------------
    assign hit_miss_set = line_hit_miss;

    //----------------------------------------------------------------------
    // MUX‐out the “data” byte from whichever way “sel” picks:
    //----------------------------------------------------------------------
    mux4to1 #(
        .w(8)
    ) mux_data_inst (
        .in_0(line_data[7:0]),
        .in_1(line_data[15:8]),
        .in_2(line_data[23:16]),
        .in_3(line_data[31:24]),
        .sel (sel),
        .out (data)
    );

    //----------------------------------------------------------------------
    // MUX‐out the “hit_miss” bit from whichever way “sel” picks:
    //----------------------------------------------------------------------
    mux4to1 #(
        .w(1)
    ) mux_hitmiss_inst (
        .in_0(line_hit_miss[0]),
        .in_1(line_hit_miss[1]),
        .in_2(line_hit_miss[2]),
        .in_3(line_hit_miss[3]),
        .sel (sel),
        .out (hit_miss)
    );

    //----------------------------------------------------------------------
    // Single clocked block for “ready” with asynchronous active‐low reset:
    //----------------------------------------------------------------------
    always @(posedge clk or negedge rst_b) begin
        if (!rst_b) begin
            // On reset, no way is “ready” to be accessed
            ready <= 4'b0000;
        end else begin
            // 1) If any way is a hit⇨ pick that way immediately (priority 0→3)
            if (line_hit_miss[0]) ready <= 4'b0001;
            else if (line_hit_miss[1]) ready <= 4'b0010;
            else if (line_hit_miss[2]) ready <= 4'b0100;
            else if (line_hit_miss[3]) ready <= 4'b1000;
            // 2) Else if no hit, pick the first empty line you find (0→3)
            else if (line_is_empty[0]) ready <= 4'b0001;
            else if (line_is_empty[1]) ready <= 4'b0010;
            else if (line_is_empty[2]) ready <= 4'b0100;
            else if (line_is_empty[3]) ready <= 4'b1000;
            // 3) Else if no empties, pick the LRU line by inspecting “ages”
            else if (ages[1:0] == 2'b11) ready <= 4'b0001;  // way0 is LRU
            else if (ages[3:2] == 2'b11) ready <= 4'b0010;  // way1 is LRU
            else if (ages[5:4] == 2'b11) ready <= 4'b0100;  // way2 is LRU
            else if (ages[7:6] == 2'b11) ready <= 4'b1000;  // way3 is LRU
            // 4) Otherwise, no line is selected (stall?)
            else
                ready <= 4'b0000;
        end
    end

endmodule
